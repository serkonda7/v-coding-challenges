module paranoia

fn test_get_inconsistencies() {
}
